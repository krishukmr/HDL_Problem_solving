//Create a module that implements a NOR gate
module top_module( 
    input a, 
    input b, 
    output out );
    nor (out,a,b);

endmodule